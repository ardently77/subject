module seg(
	input wire[3:0]a,
	output reg[6:0]b
);
  always@(*)begin
		case(a)
			4'b0000:b=7'b1000000;
			4'b0001:b=7'b1111001;
			4'b0010:b=7'b0100100;
			4'b0011:b=7'b0110000;
			4'b0100:b=7'b0011001;
			4'b0101:b=7'b0010010;
			4'b0110:b=7'b0000010;
			4'b0111:b=7'b1111000;
			4'b1000:b=7'b0000000;
			4'b1001:b=7'b0010000;
			4'b1010:b=7'b0001000;
			4'b1011:b=7'b0000011;
			4'b1100:b=7'b1000110;
			4'b1101:b=7'b0100001;
			4'b1110:b=7'b0000110;
			4'b1111:b=7'b0001110;
			default:b=7'b1000000;
		endcase
	end
endmodule
